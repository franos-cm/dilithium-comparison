`timescale 1ns / 1ps

module tb_keygen;
    localparam HIGH_PERF = 0;
    localparam SEC_LEVEL = 5;
    localparam MODE = 0;
    localparam NUM_TV = 1;

    localparam P = 10;
    localparam W = (HIGH_PERF) ? 64 : 32;

    localparam S1_SIZE = (SEC_LEVEL == 2) ? 3072
                        : (SEC_LEVEL == 3 ? 5120 : 5376);
    localparam S2_SIZE = (SEC_LEVEL == 2) ? 3072
                        : (SEC_LEVEL == 3 ? 6144 : 6144);
    localparam T0_SIZE = (SEC_LEVEL == 2) ? 13312
                        : (SEC_LEVEL == 3 ? 19968 : 26624);
    localparam T1_SIZE = (SEC_LEVEL == 2) ? 10240
                        : (SEC_LEVEL == 3 ? 15360 : 20480);
    // Ceil division for words
    localparam S1_WORDS_NUM = (S1_SIZE + W - 1) / W;
    localparam S2_WORDS_NUM = (S2_SIZE + W - 1) / W;
    localparam T0_WORDS_NUM = (T0_SIZE + W - 1) / W;
    localparam T1_WORDS_NUM = (T1_SIZE + W - 1) / W;
    localparam SEED_WORDS_NUM = (256 + W - 1) / W;
  
    logic [0:255] seed        [NUM_TV-1:0];
    logic [0:255] k           [NUM_TV-1:0];
    logic [0:255] rho         [NUM_TV-1:0];
    logic [0:255] tr          [NUM_TV-1:0];
    logic [0:S1_SIZE-1] s1    [NUM_TV-1:0];
    logic [0:S2_SIZE-1] s2    [NUM_TV-1:0];
    logic [0:T0_SIZE-1] t0    [NUM_TV-1:0];
    logic [0:T1_SIZE-1] t1    [NUM_TV-1:0];

    logic tb_rst;
    logic [9:0] ctr, c;
    integer start_time, dump_time;
    logic low_res_sk_done;

    logic clk = 1;
    logic [1:0] mode = MODE;
    logic rst, start, done;
    logic valid_i,  ready_o;
    logic ready_i, valid_o;
    logic  [W-1:0] data_i;  
    logic [W-1:0] data_o;
  
    // NOTE: different Dilithiums will have different transitions
    typedef enum logic [3:0] {
        S_INIT, S_START, S_Z, S_RHO, S_K,
        S_S1, S_S2, S_T1, S_T0, S_TR, S_STOP
    } state_t;
    state_t state;


    dilithium #(
        .HIGH_PERF(HIGH_PERF),
        .SEC_LEVEL(SEC_LEVEL)
    )
    dut (
        .clk (clk),
        .rst (rst),
        .start (start),
        .mode (mode),
        .valid_i (valid_i),
        .ready_i (ready_i),
        .data_i (data_i),
        .valid_o (valid_o),
        .ready_o (ready_o),
        .data_o (data_o)
    );
  
    initial begin
        $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/shared/seed.txt", seed);
        $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/shared/k.txt", k);
        $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/shared/rho.txt", rho);
        if (SEC_LEVEL == 2) begin
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/s1_2.txt",  s1);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/s2_2.txt",  s2);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/t0_2.txt",   t0);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/t1_2.txt",  t1);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/tr_2.txt",  tr);
        end
        else if (SEC_LEVEL == 3) begin
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/s1_3.txt",  s1);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/s2_3.txt",  s2);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/t0_3.txt",   t0);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/t1_3.txt",  t1);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/tr_3.txt",  tr);
        end
        else begin
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/s1_5.txt",  s1);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/s2_5.txt",  s2);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/t0_5.txt",   t0);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/t1_5.txt",  t1);
            $readmemh("/home/franos/projects/dilithium-comparison/tb/KAT/tr_5.txt",  tr);
        end
    end

    initial begin
        tb_rst = 1;
        #(2*P);
        tb_rst = 0;
    end

    always_ff @(posedge clk) begin
        if (tb_rst) begin
            valid_i         <= 0;
            ready_o         <= 0;
            data_i          <= 0;
            ctr             <= 0; 
            c               <= 0;
            start           <= 0;
            low_res_sk_done <= 0;
            rst             <= 1;
            state           <= S_INIT;
        end

        else begin
            rst     <= 0;
            start   <= 0;
            valid_i <= 0;
            ready_o <= 0;
            data_i  <= 0;
        
            unique case (state)
                S_INIT: begin
                    rst <= 1;
                    ctr <= ctr + 1;
                    // Arbitrary number of reset cycles
                    if (ctr == 3) begin
                        ctr <= 0;
                        state <= S_START;
                    end
                end
                S_START: begin
                    start_time <= $time;
                    start <= 1;
                    state <= S_Z;
                end
                S_Z: begin
                    valid_i <= 1;
                    data_i  <= seed[c][0 +: W];
                
                    if (ready_i) begin
                        ctr <= ctr + 1;
                        data_i <= seed[c][(ctr+1)*W +: W];

                        if (ctr == SEED_WORDS_NUM - 1) begin
                            ctr <= 0;
                            state <= S_RHO;
                        end
                    end
                end
                S_RHO: begin
                    ready_o <= 1;
                    if (valid_o) begin
                        // Since low-res dilithium dumps the data as a separate operation
                        // it is usful to keep track of both also separately
                        dump_time  <= $time;

                        if (data_o !== rho[c][ctr*W+:W])
                            $display("[Rho, %d] Error: Expected %h, received %h", ctr, rho[c][ctr*W+:W], data_o); 
                    
                        ctr <= ctr + 1;
                        
                        if (ctr == SEED_WORDS_NUM-1) begin
                            ctr <= 0;
                            state <= low_res_sk_done ? S_T1 : S_K;
                            low_res_sk_done <= !(HIGH_PERF);
                        end
                    end
                end        
                S_K: begin
                    ready_o <= 1;
                    if (valid_o) begin
                        if (data_o !== k[c][ctr*W+:W])
                            $display("[K, %d] Error: Expected %h, received %h", ctr, k[c][ctr*W+:W], data_o); 
                    
                        ctr <= ctr + 1;
                        
                        if (ctr == SEED_WORDS_NUM-1) begin
                            ctr <= 0;
                            state <= HIGH_PERF ? S_S1 : S_TR;
                        end
                    end
                end
                S_S1: begin
                    ready_o <= 1;
                    if (valid_o) begin
                        if (data_o !== s1[c][ctr*W+:W])
                            $display("[S1, %d] Error: Expected %h, received %h", ctr, s1[c][ctr*W+:W], data_o); 
        
                        ctr <= ctr + 1;
                        
                        if (ctr == S1_WORDS_NUM-1) begin
                            ctr <= 0;
                            state <= S_S2;
                        end
                    end
                end
                S_S2: begin
                    ready_o <= 1;
                    if (valid_o) begin
                        if (data_o !== s2[c][ctr*W+:W])
                            $display("[S2, %d] Error: Expected %h, received %h", ctr, s2[c][ctr*W+:W], data_o); 
                    
                        ctr <= ctr + 1;
                        
                        if (ctr == S2_WORDS_NUM-1) begin
                            ctr <= 0;
                            state <= HIGH_PERF ? S_T1 : S_T0; // S_STOP
                        end
                    end
                end
                S_T1: begin
                    ready_o <= 1;
                    if (valid_o) begin
                        if (data_o !== t1[c][ctr*W+:W])
                            $display("[T1, %d] Error: Expected %h, received %h", ctr, t1[c][ctr*W+:W], data_o); 

                        ctr <= ctr + 1;
                        
                        if (ctr == T1_WORDS_NUM-1) begin
                            ctr <= 0;
                            state <= HIGH_PERF ? S_T0 : S_STOP;
                        end
                    end
                end
                S_T0: begin
                    ready_o <= 1;
                    if (valid_o) begin
                        if (data_o !== t0[c][ctr*W+:W])
                            $display("[T0, %d] Error: Expected %h, received %h", ctr, t0[c][ctr*W+:W], data_o); 
                        ctr <= ctr + 1;
                        
                        if (ctr == T0_WORDS_NUM-1) begin
                            ctr <= 0;
                            state <= HIGH_PERF ? S_TR : S_RHO;
                        end
                    end
                end
                S_TR: begin
                    ready_o <= 1;
                    if (valid_o) begin
                        if (data_o !== tr[c][ctr*W+:W])
                            $display("[TR, %d] Error: Expected %h, received %h", ctr, tr[c][ctr*W+:W], data_o); 
                    
                        ctr <= ctr + 1;
                        
                        if (ctr == SEED_WORDS_NUM-1) begin
                            ctr <= 0;
                            state <= HIGH_PERF ? S_STOP : S_S1;
                        end
                    end
                end
                S_STOP: begin
                    ready_o <= 1;
                    c       <= c + 1;
                    state   <= S_INIT;

                    if (HIGH_PERF) begin
                        $display("KG%d[%d] completed in %d clock cycles", SEC_LEVEL, c, ($time-start_time)/P);
                    end else begin
                        $display(
                            "KG%d[%d] completed in %d (exec) + %d (dump) = %d (total) clock cycles",
                            SEC_LEVEL, c, (dump_time-start_time)/P, ($time-dump_time)/P, ($time-start_time)/P
                        );
                    end

                    if (c == NUM_TV-1) begin
                        $display ("Testbench done!");
                        $finish;
                    end
                end
                default: begin
                    $fatal(1, "Invalid state reached: %0d", state);
                end
            endcase
        end
    end
      
  
    always #(P/2) clk = ~clk;
  

endmodule