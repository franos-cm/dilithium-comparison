-- COPYRIGHT (c) 2021 ALL RIGHT RESERVED
-- Chair for Security Engineering
-- Georg Land (georg.land@rub.de)
-- License: see LICENSE file

-- THIS CODE AND INFORMATION ARE PROVIDED "AS IS" WITHOUT WARRANTY OF ANY 
-- KIND, EITHER EXPRESSED OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND/OR FITNESS FOR A
-- PARTICULAR PURPOSE.

LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.NUMERIC_STD.ALL;
LIBRARY UNISIM;
    USE UNISIM.vcomponents.ALL;
LIBRARY UNIMACRO;
    USE unimacro.Vcomponents.ALL;
    
library work;
use work.dilithium_v.all;
use work.interfaces_v.all;

entity mem_twiddle_v is
    port (
        clk : in std_logic;
        d   : in mem_twiddle_in_type;
        q   : out mem_twiddle_out_type
    );
end mem_twiddle_v;

architecture Behavioral of mem_twiddle_v is

    type tmpout_type is array(0 to 1) of std_logic_vector(31 downto 0);
    signal tmpout : tmpout_type;
    type tmpinaddr_type is array(0 to 1) of std_logic_vector(15 downto 0);
    signal tmpinaddr : tmpinaddr_type;
    
    type omegas_type is array(0 to 511) of std_logic_vector(22 downto 0);
    constant omegas : omegas_type := (
"10010010101111000000010",
"01110010111010101100111",
"01110010110010101101001",
"10011110000011000101011",
"10011111110000000110011",
"10100111101111101110011",
"10011110000011001101011",
"11101101011000110101110",
"01110010111001010000011",
"01010001110110110110000",
"00010001000000110010010",
"01101100000110111010101",
"11100001000100101001010",
"01000000111111111100100",
"11011010011110111001000",
"10011000111001010010100",
"10011101001111100011101",
"10010100001100010100111",
"11101100001000110111101",
"01010001010001111010010",
"01001010111000111011111",
"00010100101001011101110",
"01010101111011010010111",
"10000011110000010110100",
"00110100010100001110111",
"11110010100000000110100",
"10010010010101110110111",
"11001100101001010001010",
"00101100100100111101110",
"11010110111110110000001",
"01000101101100011010101",
"01101101111011100101010",
"01101000001110000011101",
"00001100000001110100100",
"10100111010101001011111",
"10100000110100001011111",
"01110010101001011110110",
"00111111001110100010101",
"01011001000001111011010",
"01010011101000100111111",
"11100110110011010000001",
"00100001011011100101100",
"00010000111111100111000",
"01110001000011111110111",
"11001011010110100000101",
"01100010111011111110100",
"01100110000111000101011",
"01100001001000100011110",
"00110101101100001110011",
"00011100010101111101101",
"01100001011011000100010",
"01000000001000010100010",
"11000100101011001001010",
"10000101000110011010100",
"00111000100100101101110",
"10010010010011001110011",
"10010010101010100111111",
"10010100101111100110101",
"01110110000111001101101",
"00100011011001011000011",
"10000111001101000011100",
"01000001110011000010010",
"00111000101101101110000",
"01011101110001111110001",
"10110001000010011001100",
"00101110101000100000010",
"00101001011001010100000",
"01001100100100010110100",
"11010111100010011010011",
"10000000100110011101000",
"00001010101001010001100",
"01111111101010101001100",
"01101010010001001011110",
"11101110011111010011110",
"10010101111011001110000",
"01010101110010110011011",
"01110111000100000100000",
"00110100111111001111001",
"10001011001101101111110",
"10101111010100100110000",
"10110110110001111010000",
"00100011000011110111010",
"01010001111000110000110",
"00111011001000010100010",
"01011100101001101001100",
"00111100101010011100110",
"00011110110111000010111",
"10100000011111011100001",
"11011000000100111010001",
"01001011001001011101100",
"11101011110100000100110",
"11011101111000111110101",
"01011001010010011111000",
"10011100100100000010111",
"10111011011111011001011",
"00100110111111010111001",
"00110110100100000100111",
"00001110101110101011001",
"10101011000010100110110",
"00111101111001001010110",
"01001011000111011001011",
"10010101010010110000010",
"11110101101111101011001",
"10011101011001011101010",
"10000000000110001111110",
"00000101001011011011000",
"01000110100101010000110",
"10100100101100010011100",
"11011010010100001011100",
"00000111001011110001111",
"11000101000101100110100",
"01110101100011011101111",
"10111010111100001111010",
"10100101010110010101001",
"10101010111100101011101",
"10001011010011011010100",
"00010010111101001101100",
"10011110001011011000001",
"10110111111001111011010",
"11110111011000101110101",
"10110111101010100110010",
"10011001111111100010010",
"11110001101111001100110",
"01111110111001010001000",
"01100110111110010101010",
"01100011011100001011001",
"00110101001111001111011",
"00000000000011011011001",
"11001110001101011000111",
"10000001001101110101001",
"01111001111010000101111",
"11111110111001101011101",
"10100011001010101110011",
"01011011011111111001011",
"10111101000100010000101",
"00100100000101000100011",
"11010010101011010001000",
"01110010010110110110010",
"01011110110001100010110",
"11001100010100101100000",
"01111001011110100110111",
"11110001110000000001101",
"11110110100000001100100",
"01010001001100000111000",
"00010001111001000000001",
"01001000110111000111001",
"01100110101001011010110",
"11000011010101110011000",
"10110000000000110001100",
"11010110011001101110101",
"10100011110000011101101",
"10000110111111111111000",
"00001111100000000010111",
"01100001100001100011100",
"00011010001111111110000",
"10010011011000011100011",
"00110010110100100100110",
"00111110001110101101000",
"00111001111111000010100",
"10101110100101100111100",
"10110111010010011111111",
"01000010111011000101010",
"11010101111011001101100",
"00011110110011011010101",
"01010000110011110111010",
"11111101000001100101100",
"01000111111110001100101",
"00010011011011111111111",
"01001100000001110111101",
"00100101110101101100111",
"00001111100000011110001",
"01010001101111000000110",
"11001110011100101010111",
"01111011010011000000100",
"10000110011101010101100",
"11111101111100011110101",
"00010000000111001101101",
"11110111100011101011001",
"00010000101001001100000",
"10000110111111100110001",
"00010110111000000001001",
"11010111110000111001100",
"01011001010010111100110",
"10011011100000001001110",
"11101001101000010111101",
"00100110010001100101110",
"00000100010001111010100",
"11111000000110110110011",
"00100011100000101001110",
"11100110110000110111000",
"00100000001011100001110",
"11000100101011111000101",
"01000000001111111000110",
"11001001101001111010101",
"11111111011000110011010",
"00011001000110100001101",
"11110101011011000001101",
"00000100010101000001011",
"01011111010101000110010",
"00000010101010010101000",
"00111100110110100111110",
"01000110000100100100011",
"11011110000101000010001",
"10010111101010101111001",
"01001110011001100110011",
"11000101000110000110111",
"01101011110000111011101",
"11001001011010111111110",
"11011011110000000100100",
"10010001100001110011011",
"00000110100011101100000",
"00110000101110110010110",
"01111110100110011110101",
"00010010101101101110110",
"11001011010110110110011",
"10111001101010110110100",
"11011011011111111010100",
"01010000101010000100100",
"01101000101100000100100",
"00010011011010000110100",
"00111101111001000000110",
"11000110011000010111011",
"11100111111000111001110",
"11010011010100011101111",
"11000001101011101110010",
"11001011000010110010001",
"01011100001011001101001",
"10110100110110110000000",
"01011011110110011010100",
"01001100101100001111010",
"10111100110100101000010",
"10000110101111010000111",
"11010101001110111111010",
"10001010100110111110010",
"11101110110110100001011",
"10001100101110110001101",
"00110100100101101011101",
"10010101110010100111100",
"10001100100101011011110",
"01010100100111001111000",
"10101100000001110001110",
"10011110101100001011001",
"11101000001111001111000",
"10001101000001010011000",
"10000100111111000100011",
"10111100000011000011110",
"11110011110000111111110",
"10001110010100010101111",
"11000111110000111100011",
"11111111010111110000000",
"11010001100010101011001",
"10110100110100010110000",
"10011000111011011001000",
"10111101010000001101100",
"11101001011011011010111",
"00000000000000000000000",
"00001011001010010010101",
"10100001000111111001011",
"10110011010010010011101",
"10100101010101110101001",
"00010111000110101010100",
"10000000000100001000001",
"00011011111111100001111",
"00111000101101110101001",
"10000101110111100000010",
"10100001101110011110010",
"00111101011000011101111",
"10111001001111010110101",
"10001011101000011000101",
"00110000100001111010100",
"10101001101111000111010",
"11010101011100011000101",
"10111001011101010010010",
"10110100110110101100011",
"01100101100101001010010",
"00111001100000100111010",
"00001000011100101111011",
"10111010011100100001000",
"10010101001000100000100",
"00111100100000010111101",
"10100001010101101100000",
"11011001011001111000100",
"11010001110100110010111",
"10100101010100101000001",
"01010001110010011001100",
"00011010010110100111000",
"10011110111010001001000",
"00010110001101110001001",
"10001011110011100011010",
"00011100101011110100011",
"11100000110011011111110",
"11110110000010111100111",
"11001011011001111101111",
"11010111011010111101111",
"10010010000000000010111",
"10100010111010100100111",
"00011010001100100100111",
"11110110011001001000110",
"01000000100100110000110",
"11100111011000100110110",
"11111100011110001010001",
"00110111000111000110011",
"10010001110111111101111",
"10011011000010100000010",
"01001001111111100010010",
"00011101010100111100101",
"01011000101011001100111",
"00110100000010101000100",
"00010000110101011111000",
"01011100110101101101111",
"11100001010100101100010",
"11111110011010110101101",
"11010000000101011101000",
"01111101101101011111011",
"00000101001010011111010",
"01110011010100101111010",
"10000000000011100110100",
"00011011000011000010110",
"11011111101000000011110",
"00011101100010000011110",
"11101111101010001111010",
"10001100010111100100101",
"11101101111111101011010",
"00000011110100100100111",
"11111101100111000010111",
"11101100100111001101010",
"00001011000011110100010",
"10110001111111111011010",
"11010011000110100001110",
"10010011110111100011011",
"01110100011011111111100",
"00111100011000001101000",
"11110111011011011010001",
"00000100000110001010100",
"01110111110100011001010",
"00000000111001110000110",
"10111100100001010101011",
"11000010000110011111111",
"00011000101001101010101",
"11010110111000011111110",
"01111000000111110001000",
"01101100111101001001101",
"01011001110111000100010",
"01110110001010000000001",
"01011011111000111001110",
"10000001001111001101011",
"11010111010110000100100",
"01110000011110010010110",
"10010100110010011001011",
"11011110010010011101100",
"00100100001110110000001",
"10101000011101001100011",
"11100010110000011110111",
"11100000101000101001101",
"11100110010101101101110",
"00110110001011110001111",
"11110010101000000001001",
"11001110111111001110011",
"01111000000111111110101",
"10111100010000000000101",
"00101101111111110001010",
"00010100101011001000110",
"10100111101111100111011",
"10011110000101000110101",
"11001100011011010010110",
"01011011011100011100100",
"01110110111011100000000",
"11010111001001111100101",
"10000100011111111001111",
"00000110111111111111010",
"01000011001000101100101",
"10011001100101101010001",
"11010000010111001110110",
"11000110100100100101000",
"10010110011010010111101",
"01101101110101011101111",
"00100001010101110111110",
"01010010001000000011011",
"00101110010010101000111",
"00000000011011001010010",
"01000010111010111101001",
"00111111010001000101100",
"00011000110001010011101",
"01111111110110010010100",
"01100101010000011000011",
"01001110001001111010100",
"11001100010000110101100",
"11000000010011010111101",
"10000110111000011001110",
"10110010110000001111000",
"10100011111010101101000",
"00000100001011101000110",
"10100011110011000010100",
"00110000110010010100000",
"11110110010001011001011",
"10111010000110010010111",
"00101010011001101010010",
"00101101001100110101100",
"10100010010001111000100",
"01000101000110010001001",
"10011101001101001100111",
"01111100010010000111001",
"10010010100101111010011",
"10101101011001110110011",
"11011100011101010111110",
"11111101001010010010101",
"10111111101100111000010",
"10110001000011010001100",
"00000101000000001010100",
"10110101000110101000000",
"01011010010100010011011",
"11100000110011011010110",
"10101010001110101100110",
"01111000100000101010100",
"01100100100101111101101",
"01101100011000010100100",
"00100010001000010011011",
"00110001100101111110101",
"11010011000110110000101",
"00010000111011100000110",
"10001001110101111101110",
"11011010001011010001011",
"00010011110101100011000",
"00101111101000010010000",
"01110000011100011110101",
"11100001011010110001110",
"11010001011011001011011",
"11100010001011110110000",
"11010110110011100111110",
"11101110001110000100100",
"10100100010111000011001",
"10101000000101101101001",
"10111010001001001000010",
"01100101011000011000100",
"11000100001101111110001",
"01010100111110100110011",
"10110100110010011001001",
"10001000100000010110010",
"11001010100111011010010",
"10111111111010101011011",
"11111010011011010111011",
"10111111011100110001101",
"00010100000110110010111",
"11011001011101110100111",
"11101011000011010110001",
"11101000011011110000000",
"10100111001110110011011",
"01010000111111000001000",
"11100011011001001001001",
"11011110110110011111000",
"10111100001001011110011",
"01101110001011010011111",
"01000100110100011001010",
"00110101100000001100110",
"00110110100010101100001",
"00110110101110011000111",
"11100011011101101001010",
"10111101001100110010111",
"10011101011010011011100",
"11011111101011110110000",
"11001111000010011110000",
"01110001101101000001010",
"01100101000001111000111",
"11001111001011101110010",
"01001100110100011101011",
"11001110010010000000111",
"00011010001100101111110",
"01000111010110000000101",
"11110111010000001100101",
"11101111000010001101011",
"00001100011110011000000",
"01010110000011101100001",
"11010011001111000010100",
"01100000010000101110110",
"11000110011011010000110",
"00101111011101111010001",
"00101100001101011010001",
"11111001101111000101111",
"01001011110000111110010",
"11001000110010001101100",
"01011101000001110010110",
"00010100011000101000000",
"11101001011101100001010",
"10011001011011010111100",
"00110110101101000100101",
"10000110011111111100111",
"01100101101101111000101",
"10111101110111110100111",
"01010100111010010110101",
"11110101011011010001010",
"01011010011011100010001",
"11010111000111000011000",
"00001001110011100100010",
"00110101110001110101101",
"00110001010000001110010",
"10110011010011010110111",
"10010010100000100011101",
"11011111010000000001111",
"10001111001101101011100",
"01001001110100100010110",
"11110111001111100111000",
"11010110110100100101001",
"01000110011011010111111",
"10001001000011100101010",
"00110000110110011001011",
"00101100000000001000111",
"00101111111111111100111",
"00110000110110011101011",
"01000110011110101001100",
"01000110011010101001101",
"10110110011000100000000",
"00000000000000000000000"
);

    type init_type is array(0 to 63) of std_logic_vector(255 downto 0);
    constant init : init_type := (
"000000000" & omegas(7) & "000000000" & omegas(6) & "000000000" & omegas(5) & "000000000" & omegas(4) & "000000000" & omegas(3) & "000000000" & omegas(2) & "000000000" & omegas(1) & "000000000" & omegas(0),
"000000000" & omegas(15) & "000000000" & omegas(14) & "000000000" & omegas(13) & "000000000" & omegas(12) & "000000000" & omegas(11) & "000000000" & omegas(10) & "000000000" & omegas(9) & "000000000" & omegas(8),
"000000000" & omegas(23) & "000000000" & omegas(22) & "000000000" & omegas(21) & "000000000" & omegas(20) & "000000000" & omegas(19) & "000000000" & omegas(18) & "000000000" & omegas(17) & "000000000" & omegas(16),
"000000000" & omegas(31) & "000000000" & omegas(30) & "000000000" & omegas(29) & "000000000" & omegas(28) & "000000000" & omegas(27) & "000000000" & omegas(26) & "000000000" & omegas(25) & "000000000" & omegas(24),
"000000000" & omegas(39) & "000000000" & omegas(38) & "000000000" & omegas(37) & "000000000" & omegas(36) & "000000000" & omegas(35) & "000000000" & omegas(34) & "000000000" & omegas(33) & "000000000" & omegas(32),
"000000000" & omegas(47) & "000000000" & omegas(46) & "000000000" & omegas(45) & "000000000" & omegas(44) & "000000000" & omegas(43) & "000000000" & omegas(42) & "000000000" & omegas(41) & "000000000" & omegas(40),
"000000000" & omegas(55) & "000000000" & omegas(54) & "000000000" & omegas(53) & "000000000" & omegas(52) & "000000000" & omegas(51) & "000000000" & omegas(50) & "000000000" & omegas(49) & "000000000" & omegas(48),
"000000000" & omegas(63) & "000000000" & omegas(62) & "000000000" & omegas(61) & "000000000" & omegas(60) & "000000000" & omegas(59) & "000000000" & omegas(58) & "000000000" & omegas(57) & "000000000" & omegas(56),
"000000000" & omegas(71) & "000000000" & omegas(70) & "000000000" & omegas(69) & "000000000" & omegas(68) & "000000000" & omegas(67) & "000000000" & omegas(66) & "000000000" & omegas(65) & "000000000" & omegas(64),
"000000000" & omegas(79) & "000000000" & omegas(78) & "000000000" & omegas(77) & "000000000" & omegas(76) & "000000000" & omegas(75) & "000000000" & omegas(74) & "000000000" & omegas(73) & "000000000" & omegas(72),
"000000000" & omegas(87) & "000000000" & omegas(86) & "000000000" & omegas(85) & "000000000" & omegas(84) & "000000000" & omegas(83) & "000000000" & omegas(82) & "000000000" & omegas(81) & "000000000" & omegas(80),
"000000000" & omegas(95) & "000000000" & omegas(94) & "000000000" & omegas(93) & "000000000" & omegas(92) & "000000000" & omegas(91) & "000000000" & omegas(90) & "000000000" & omegas(89) & "000000000" & omegas(88),
"000000000" & omegas(103) & "000000000" & omegas(102) & "000000000" & omegas(101) & "000000000" & omegas(100) & "000000000" & omegas(99) & "000000000" & omegas(98) & "000000000" & omegas(97) & "000000000" & omegas(96),
"000000000" & omegas(111) & "000000000" & omegas(110) & "000000000" & omegas(109) & "000000000" & omegas(108) & "000000000" & omegas(107) & "000000000" & omegas(106) & "000000000" & omegas(105) & "000000000" & omegas(104),
"000000000" & omegas(119) & "000000000" & omegas(118) & "000000000" & omegas(117) & "000000000" & omegas(116) & "000000000" & omegas(115) & "000000000" & omegas(114) & "000000000" & omegas(113) & "000000000" & omegas(112),
"000000000" & omegas(127) & "000000000" & omegas(126) & "000000000" & omegas(125) & "000000000" & omegas(124) & "000000000" & omegas(123) & "000000000" & omegas(122) & "000000000" & omegas(121) & "000000000" & omegas(120),
"000000000" & omegas(135) & "000000000" & omegas(134) & "000000000" & omegas(133) & "000000000" & omegas(132) & "000000000" & omegas(131) & "000000000" & omegas(130) & "000000000" & omegas(129) & "000000000" & omegas(128),
"000000000" & omegas(143) & "000000000" & omegas(142) & "000000000" & omegas(141) & "000000000" & omegas(140) & "000000000" & omegas(139) & "000000000" & omegas(138) & "000000000" & omegas(137) & "000000000" & omegas(136),
"000000000" & omegas(151) & "000000000" & omegas(150) & "000000000" & omegas(149) & "000000000" & omegas(148) & "000000000" & omegas(147) & "000000000" & omegas(146) & "000000000" & omegas(145) & "000000000" & omegas(144),
"000000000" & omegas(159) & "000000000" & omegas(158) & "000000000" & omegas(157) & "000000000" & omegas(156) & "000000000" & omegas(155) & "000000000" & omegas(154) & "000000000" & omegas(153) & "000000000" & omegas(152),
"000000000" & omegas(167) & "000000000" & omegas(166) & "000000000" & omegas(165) & "000000000" & omegas(164) & "000000000" & omegas(163) & "000000000" & omegas(162) & "000000000" & omegas(161) & "000000000" & omegas(160),
"000000000" & omegas(175) & "000000000" & omegas(174) & "000000000" & omegas(173) & "000000000" & omegas(172) & "000000000" & omegas(171) & "000000000" & omegas(170) & "000000000" & omegas(169) & "000000000" & omegas(168),
"000000000" & omegas(183) & "000000000" & omegas(182) & "000000000" & omegas(181) & "000000000" & omegas(180) & "000000000" & omegas(179) & "000000000" & omegas(178) & "000000000" & omegas(177) & "000000000" & omegas(176),
"000000000" & omegas(191) & "000000000" & omegas(190) & "000000000" & omegas(189) & "000000000" & omegas(188) & "000000000" & omegas(187) & "000000000" & omegas(186) & "000000000" & omegas(185) & "000000000" & omegas(184),
"000000000" & omegas(199) & "000000000" & omegas(198) & "000000000" & omegas(197) & "000000000" & omegas(196) & "000000000" & omegas(195) & "000000000" & omegas(194) & "000000000" & omegas(193) & "000000000" & omegas(192),
"000000000" & omegas(207) & "000000000" & omegas(206) & "000000000" & omegas(205) & "000000000" & omegas(204) & "000000000" & omegas(203) & "000000000" & omegas(202) & "000000000" & omegas(201) & "000000000" & omegas(200),
"000000000" & omegas(215) & "000000000" & omegas(214) & "000000000" & omegas(213) & "000000000" & omegas(212) & "000000000" & omegas(211) & "000000000" & omegas(210) & "000000000" & omegas(209) & "000000000" & omegas(208),
"000000000" & omegas(223) & "000000000" & omegas(222) & "000000000" & omegas(221) & "000000000" & omegas(220) & "000000000" & omegas(219) & "000000000" & omegas(218) & "000000000" & omegas(217) & "000000000" & omegas(216),
"000000000" & omegas(231) & "000000000" & omegas(230) & "000000000" & omegas(229) & "000000000" & omegas(228) & "000000000" & omegas(227) & "000000000" & omegas(226) & "000000000" & omegas(225) & "000000000" & omegas(224),
"000000000" & omegas(239) & "000000000" & omegas(238) & "000000000" & omegas(237) & "000000000" & omegas(236) & "000000000" & omegas(235) & "000000000" & omegas(234) & "000000000" & omegas(233) & "000000000" & omegas(232),
"000000000" & omegas(247) & "000000000" & omegas(246) & "000000000" & omegas(245) & "000000000" & omegas(244) & "000000000" & omegas(243) & "000000000" & omegas(242) & "000000000" & omegas(241) & "000000000" & omegas(240),
"000000000" & omegas(255) & "000000000" & omegas(254) & "000000000" & omegas(253) & "000000000" & omegas(252) & "000000000" & omegas(251) & "000000000" & omegas(250) & "000000000" & omegas(249) & "000000000" & omegas(248),
"000000000" & omegas(263) & "000000000" & omegas(262) & "000000000" & omegas(261) & "000000000" & omegas(260) & "000000000" & omegas(259) & "000000000" & omegas(258) & "000000000" & omegas(257) & "000000000" & omegas(256),
"000000000" & omegas(271) & "000000000" & omegas(270) & "000000000" & omegas(269) & "000000000" & omegas(268) & "000000000" & omegas(267) & "000000000" & omegas(266) & "000000000" & omegas(265) & "000000000" & omegas(264),
"000000000" & omegas(279) & "000000000" & omegas(278) & "000000000" & omegas(277) & "000000000" & omegas(276) & "000000000" & omegas(275) & "000000000" & omegas(274) & "000000000" & omegas(273) & "000000000" & omegas(272),
"000000000" & omegas(287) & "000000000" & omegas(286) & "000000000" & omegas(285) & "000000000" & omegas(284) & "000000000" & omegas(283) & "000000000" & omegas(282) & "000000000" & omegas(281) & "000000000" & omegas(280),
"000000000" & omegas(295) & "000000000" & omegas(294) & "000000000" & omegas(293) & "000000000" & omegas(292) & "000000000" & omegas(291) & "000000000" & omegas(290) & "000000000" & omegas(289) & "000000000" & omegas(288),
"000000000" & omegas(303) & "000000000" & omegas(302) & "000000000" & omegas(301) & "000000000" & omegas(300) & "000000000" & omegas(299) & "000000000" & omegas(298) & "000000000" & omegas(297) & "000000000" & omegas(296),
"000000000" & omegas(311) & "000000000" & omegas(310) & "000000000" & omegas(309) & "000000000" & omegas(308) & "000000000" & omegas(307) & "000000000" & omegas(306) & "000000000" & omegas(305) & "000000000" & omegas(304),
"000000000" & omegas(319) & "000000000" & omegas(318) & "000000000" & omegas(317) & "000000000" & omegas(316) & "000000000" & omegas(315) & "000000000" & omegas(314) & "000000000" & omegas(313) & "000000000" & omegas(312),
"000000000" & omegas(327) & "000000000" & omegas(326) & "000000000" & omegas(325) & "000000000" & omegas(324) & "000000000" & omegas(323) & "000000000" & omegas(322) & "000000000" & omegas(321) & "000000000" & omegas(320),
"000000000" & omegas(335) & "000000000" & omegas(334) & "000000000" & omegas(333) & "000000000" & omegas(332) & "000000000" & omegas(331) & "000000000" & omegas(330) & "000000000" & omegas(329) & "000000000" & omegas(328),
"000000000" & omegas(343) & "000000000" & omegas(342) & "000000000" & omegas(341) & "000000000" & omegas(340) & "000000000" & omegas(339) & "000000000" & omegas(338) & "000000000" & omegas(337) & "000000000" & omegas(336),
"000000000" & omegas(351) & "000000000" & omegas(350) & "000000000" & omegas(349) & "000000000" & omegas(348) & "000000000" & omegas(347) & "000000000" & omegas(346) & "000000000" & omegas(345) & "000000000" & omegas(344),
"000000000" & omegas(359) & "000000000" & omegas(358) & "000000000" & omegas(357) & "000000000" & omegas(356) & "000000000" & omegas(355) & "000000000" & omegas(354) & "000000000" & omegas(353) & "000000000" & omegas(352),
"000000000" & omegas(367) & "000000000" & omegas(366) & "000000000" & omegas(365) & "000000000" & omegas(364) & "000000000" & omegas(363) & "000000000" & omegas(362) & "000000000" & omegas(361) & "000000000" & omegas(360),
"000000000" & omegas(375) & "000000000" & omegas(374) & "000000000" & omegas(373) & "000000000" & omegas(372) & "000000000" & omegas(371) & "000000000" & omegas(370) & "000000000" & omegas(369) & "000000000" & omegas(368),
"000000000" & omegas(383) & "000000000" & omegas(382) & "000000000" & omegas(381) & "000000000" & omegas(380) & "000000000" & omegas(379) & "000000000" & omegas(378) & "000000000" & omegas(377) & "000000000" & omegas(376),
"000000000" & omegas(391) & "000000000" & omegas(390) & "000000000" & omegas(389) & "000000000" & omegas(388) & "000000000" & omegas(387) & "000000000" & omegas(386) & "000000000" & omegas(385) & "000000000" & omegas(384),
"000000000" & omegas(399) & "000000000" & omegas(398) & "000000000" & omegas(397) & "000000000" & omegas(396) & "000000000" & omegas(395) & "000000000" & omegas(394) & "000000000" & omegas(393) & "000000000" & omegas(392),
"000000000" & omegas(407) & "000000000" & omegas(406) & "000000000" & omegas(405) & "000000000" & omegas(404) & "000000000" & omegas(403) & "000000000" & omegas(402) & "000000000" & omegas(401) & "000000000" & omegas(400),
"000000000" & omegas(415) & "000000000" & omegas(414) & "000000000" & omegas(413) & "000000000" & omegas(412) & "000000000" & omegas(411) & "000000000" & omegas(410) & "000000000" & omegas(409) & "000000000" & omegas(408),
"000000000" & omegas(423) & "000000000" & omegas(422) & "000000000" & omegas(421) & "000000000" & omegas(420) & "000000000" & omegas(419) & "000000000" & omegas(418) & "000000000" & omegas(417) & "000000000" & omegas(416),
"000000000" & omegas(431) & "000000000" & omegas(430) & "000000000" & omegas(429) & "000000000" & omegas(428) & "000000000" & omegas(427) & "000000000" & omegas(426) & "000000000" & omegas(425) & "000000000" & omegas(424),
"000000000" & omegas(439) & "000000000" & omegas(438) & "000000000" & omegas(437) & "000000000" & omegas(436) & "000000000" & omegas(435) & "000000000" & omegas(434) & "000000000" & omegas(433) & "000000000" & omegas(432),
"000000000" & omegas(447) & "000000000" & omegas(446) & "000000000" & omegas(445) & "000000000" & omegas(444) & "000000000" & omegas(443) & "000000000" & omegas(442) & "000000000" & omegas(441) & "000000000" & omegas(440),
"000000000" & omegas(455) & "000000000" & omegas(454) & "000000000" & omegas(453) & "000000000" & omegas(452) & "000000000" & omegas(451) & "000000000" & omegas(450) & "000000000" & omegas(449) & "000000000" & omegas(448),
"000000000" & omegas(463) & "000000000" & omegas(462) & "000000000" & omegas(461) & "000000000" & omegas(460) & "000000000" & omegas(459) & "000000000" & omegas(458) & "000000000" & omegas(457) & "000000000" & omegas(456),
"000000000" & omegas(471) & "000000000" & omegas(470) & "000000000" & omegas(469) & "000000000" & omegas(468) & "000000000" & omegas(467) & "000000000" & omegas(466) & "000000000" & omegas(465) & "000000000" & omegas(464),
"000000000" & omegas(479) & "000000000" & omegas(478) & "000000000" & omegas(477) & "000000000" & omegas(476) & "000000000" & omegas(475) & "000000000" & omegas(474) & "000000000" & omegas(473) & "000000000" & omegas(472),
"000000000" & omegas(487) & "000000000" & omegas(486) & "000000000" & omegas(485) & "000000000" & omegas(484) & "000000000" & omegas(483) & "000000000" & omegas(482) & "000000000" & omegas(481) & "000000000" & omegas(480),
"000000000" & omegas(495) & "000000000" & omegas(494) & "000000000" & omegas(493) & "000000000" & omegas(492) & "000000000" & omegas(491) & "000000000" & omegas(490) & "000000000" & omegas(489) & "000000000" & omegas(488),
"000000000" & omegas(503) & "000000000" & omegas(502) & "000000000" & omegas(501) & "000000000" & omegas(500) & "000000000" & omegas(499) & "000000000" & omegas(498) & "000000000" & omegas(497) & "000000000" & omegas(496),
"000000000" & omegas(511) & "000000000" & omegas(510) & "000000000" & omegas(509) & "000000000" & omegas(508) & "000000000" & omegas(507) & "000000000" & omegas(506) & "000000000" & omegas(505) & "000000000" & omegas(504)
);
begin

    tmpinaddr(0)(4 downto 0) <= (others => '0');
    tmpinaddr(1)(4 downto 0) <= (others => '0');
    tmpinaddr(0)(15 downto 14) <= (others => '0');
    tmpinaddr(1)(15 downto 14) <= (others => '0');
    tmpinaddr(0)(13 downto 5) <= d.addr(0);
    tmpinaddr(1)(13 downto 5) <= d.addr(1);
    q(0) <= tmpout(0)(22 downto 0);
    q(1) <= tmpout(1)(22 downto 0);

   -- RAMB36E1: 18K-bit Configurable Synchronous Block RAM
   --           Artix-7
   -- Xilinx HDL Language Template, version 2020.2

   RAMB36E1_inst : RAMB36E1
   generic map (
      -- Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
      RDADDR_COLLISION_HWCONFIG => "PERFORMANCE",
      -- Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
      SIM_COLLISION_CHECK => "ALL",
      -- DOA_REG, DOB_REG: Optional output register (0 or 1)
      DOA_REG => 0,
      DOB_REG => 0,
      EN_ECC_READ => FALSE,                                                            -- Enable ECC decoder,
                                                                                       -- FALSE, TRUE
      EN_ECC_WRITE => FALSE,                                                           -- Enable ECC encoder,
                                                                                       -- FALSE, TRUE
      -- INITP_00 to INITP_0F: Initial contents of the parity memory array
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => to_bitvector(init(0)),
        INIT_01 => to_bitvector(init(1)),
        INIT_02 => to_bitvector(init(2)),
        INIT_03 => to_bitvector(init(3)),
        INIT_04 => to_bitvector(init(4)),
        INIT_05 => to_bitvector(init(5)),
        INIT_06 => to_bitvector(init(6)),
        INIT_07 => to_bitvector(init(7)),
        INIT_08 => to_bitvector(init(8)),
        INIT_09 => to_bitvector(init(9)),
        INIT_0A => to_bitvector(init(10)),
        INIT_0B => to_bitvector(init(11)),
        INIT_0C => to_bitvector(init(12)),
        INIT_0D => to_bitvector(init(13)),
        INIT_0E => to_bitvector(init(14)),
        INIT_0F => to_bitvector(init(15)),
        INIT_10 => to_bitvector(init(16)),
        INIT_11 => to_bitvector(init(17)),
        INIT_12 => to_bitvector(init(18)),
        INIT_13 => to_bitvector(init(19)),
        INIT_14 => to_bitvector(init(20)),
        INIT_15 => to_bitvector(init(21)),
        INIT_16 => to_bitvector(init(22)),
        INIT_17 => to_bitvector(init(23)),
        INIT_18 => to_bitvector(init(24)),
        INIT_19 => to_bitvector(init(25)),
        INIT_1A => to_bitvector(init(26)),
        INIT_1B => to_bitvector(init(27)),
        INIT_1C => to_bitvector(init(28)),
        INIT_1D => to_bitvector(init(29)),
        INIT_1E => to_bitvector(init(30)),
        INIT_1F => to_bitvector(init(31)),
        INIT_20 => to_bitvector(init(32)),
        INIT_21 => to_bitvector(init(33)),
        INIT_22 => to_bitvector(init(34)),
        INIT_23 => to_bitvector(init(35)),
        INIT_24 => to_bitvector(init(36)),
        INIT_25 => to_bitvector(init(37)),
        INIT_26 => to_bitvector(init(38)),
        INIT_27 => to_bitvector(init(39)),
        INIT_28 => to_bitvector(init(40)),
        INIT_29 => to_bitvector(init(41)),
        INIT_2A => to_bitvector(init(42)),
        INIT_2B => to_bitvector(init(43)),
        INIT_2C => to_bitvector(init(44)),
        INIT_2D => to_bitvector(init(45)),
        INIT_2E => to_bitvector(init(46)),
        INIT_2F => to_bitvector(init(47)),
        INIT_30 => to_bitvector(init(48)),
        INIT_31 => to_bitvector(init(49)),
        INIT_32 => to_bitvector(init(50)),
        INIT_33 => to_bitvector(init(51)),
        INIT_34 => to_bitvector(init(52)),
        INIT_35 => to_bitvector(init(53)),
        INIT_36 => to_bitvector(init(54)),
        INIT_37 => to_bitvector(init(55)),
        INIT_38 => to_bitvector(init(56)),
        INIT_39 => to_bitvector(init(57)),
        INIT_3A => to_bitvector(init(58)),
        INIT_3B => to_bitvector(init(59)),
        INIT_3C => to_bitvector(init(60)),
        INIT_3D => to_bitvector(init(61)),
        INIT_3E => to_bitvector(init(62)),
        INIT_3F => to_bitvector(init(63)),
      INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- INIT_A, INIT_B: Initial values on output ports
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      -- Initialization File: RAM initialization file
      INIT_FILE => "NONE",
      -- RAM Mode: "SDP" or "TDP" 
      RAM_MODE => "TDP",
      -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      -- READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
      READ_WIDTH_A => 36,                                                               -- 0-72
      READ_WIDTH_B => 36,                                                               -- 0-36
      WRITE_WIDTH_A => 0,                                                              -- 0-36
      WRITE_WIDTH_B => 0,                                                              -- 0-72
      -- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
      RSTREG_PRIORITY_A => "REGCE",
      RSTREG_PRIORITY_B => "REGCE",
      -- SRVAL_A, SRVAL_B: Set/reset value for output
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      -- Simulation Device: Must be set to "7SERIES" for simulation behavior
      SIM_DEVICE => "7SERIES",
      -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
      WRITE_MODE_A => "NO_CHANGE",
      WRITE_MODE_B => "NO_CHANGE" 
   )
   port map (
      -- Cascade Signals: 1-bit (each) output: BRAM cascade ports (to create 64kx1)
      CASCADEOUTA => open,     -- 1-bit output: A port cascade
      CASCADEOUTB => open,     -- 1-bit output: B port cascade
      -- ECC Signals: 1-bit (each) output: Error Correction Circuitry ports
      DBITERR => open,             -- 1-bit output: Double bit error status
      ECCPARITY => open,         -- 8-bit output: Generated error correction parity
      RDADDRECC => open,         -- 9-bit output: ECC read address
      SBITERR => open,             -- 1-bit output: Single bit error status
      -- Port A Data: 32-bit (each) output: Port A data
      DOADO => tmpout(0),                 -- 32-bit output: A port data/LSB data
      DOPADOP => open,             -- 4-bit output: A port parity/LSB parity
      -- Port B Data: 32-bit (each) output: Port B data
      DOBDO => tmpout(1),                 -- 32-bit output: B port data/MSB data
      DOPBDOP => open,             -- 4-bit output: B port parity/MSB parity
      -- Cascade Signals: 1-bit (each) input: BRAM cascade ports (to create 64kx1)
      CASCADEINA => '0',       -- 1-bit input: A port cascade
      CASCADEINB => '0',       -- 1-bit input: B port cascade
      -- ECC Signals: 1-bit (each) input: Error Correction Circuitry ports
      INJECTDBITERR => '0', -- 1-bit input: Inject a double bit error
      INJECTSBITERR => '0', -- 1-bit input: Inject a single bit error
      -- Port A Address/Control Signals: 16-bit (each) input: Port A address and control signals (read port
      -- when RAM_MODE="SDP")
      ADDRARDADDR => tmpinaddr(0),     -- 16-bit input: A port address/Read address
      CLKARDCLK => clk,         -- 1-bit input: A port clock/Read clock
      ENARDEN => d.en(0),             -- 1-bit input: A port enable/Read enable
      REGCEAREGCE => '1',     -- 1-bit input: A port register enable/Register enable
      RSTRAMARSTRAM => '0', -- 1-bit input: A port set/reset
      RSTREGARSTREG => '0', -- 1-bit input: A port register set/reset
      WEA => (others => '0'),                     -- 4-bit input: A port write enable
      -- Port A Data: 32-bit (each) input: Port A data
      DIADI => (others => '0'),                 -- 32-bit input: A port data/LSB data
      DIPADIP => (others => '0'),             -- 4-bit input: A port parity/LSB parity
      -- Port B Address/Control Signals: 16-bit (each) input: Port B address and control signals (write port
      -- when RAM_MODE="SDP")
      ADDRBWRADDR => tmpinaddr(1),     -- 16-bit input: B port address/Write address
      CLKBWRCLK => clk,         -- 1-bit input: B port clock/Write clock
      ENBWREN => d.en(1),             -- 1-bit input: B port enable/Write enable
      REGCEB => '1',               -- 1-bit input: B port register enable
      RSTRAMB => '0',             -- 1-bit input: B port set/reset
      RSTREGB => '0',             -- 1-bit input: B port register set/reset
      WEBWE => (others => '0'),                 -- 8-bit input: B port write enable/Write enable
      -- Port B Data: 32-bit (each) input: Port B data
      DIBDI => (others => '0'),                 -- 32-bit input: B port data/MSB data
      DIPBDIP => (others => '0')              -- 4-bit input: B port parity/MSB parity
   );

   -- End of RAMB36E1_inst instantiation

end Behavioral;