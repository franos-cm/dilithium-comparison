-- COPYRIGHT (c) 2021 ALL RIGHT RESERVED
-- Chair for Security Engineering
-- Georg Land (georg.land@rub.de)
-- License: see LICENSE file

-- THIS CODE AND INFORMATION ARE PROVIDED "AS IS" WITHOUT WARRANTY OF ANY 
-- KIND, EITHER EXPRESSED OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND/OR FITNESS FOR A
-- PARTICULAR PURPOSE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
use UNISIM.VComponents.all;
Library UNIMACRO;
use UNIMACRO.vcomponents.all;

library work;
use work.dilithium_iii.all;
use work.interfaces.all;
use work.memmap_iii.all;

entity mem_8_quarter_poly is
    Port (
        clk : in std_logic;
        d   : in mem_8_quarter_poly_in_type;
        q   : out std_logic_vector(22 downto 0)
    );
end mem_8_quarter_poly;

architecture Behavioral of mem_8_quarter_poly is

--    type storage_type is array(0 to 511) of std_logic_vector(22 downto 0);
--    signal storage : storage_type := (others => (others => '0'));

--    signal din, dout : std_logic_vector(31 downto 0);
--    signal raddr, waddr : std_logic_vector(13 downto 0);

begin
--  <-----Cut code below this line and paste into the architecture body---->

   -- BRAM_SDP_MACRO: Simple Dual Port RAM
   --                 Artix-7
   -- Xilinx HDL Language Template, version 2020.1
   
   -- Note -  This Unimacro model assumes the port directions to be "downto". 
   --         Simulation of this model with "to" in the port directions could lead to erroneous results.

   -----------------------------------------------------------------------
   --  READ_WIDTH | BRAM_SIZE | READ Depth  | RDADDR Width |            --
   -- WRITE_WIDTH |           | WRITE Depth | WRADDR Width |  WE Width  --
   -- ============|===========|=============|==============|============--
   --    37-72    |  "36Kb"   |      512    |     9-bit    |    8-bit   --
   --    19-36    |  "36Kb"   |     1024    |    10-bit    |    4-bit   --
   --    19-36    |  "18Kb"   |      512    |     9-bit    |    4-bit   --
   --    10-18    |  "36Kb"   |     2048    |    11-bit    |    2-bit   --
   --    10-18    |  "18Kb"   |     1024    |    10-bit    |    2-bit   --
   --     5-9     |  "36Kb"   |     4096    |    12-bit    |    1-bit   --
   --     5-9     |  "18Kb"   |     2048    |    11-bit    |    1-bit   --
   --     3-4     |  "36Kb"   |     8192    |    13-bit    |    1-bit   --
   --     3-4     |  "18Kb"   |     4096    |    12-bit    |    1-bit   --
   --       2     |  "36Kb"   |    16384    |    14-bit    |    1-bit   --
   --       2     |  "18Kb"   |     8192    |    13-bit    |    1-bit   --
   --       1     |  "36Kb"   |    32768    |    15-bit    |    1-bit   --
   --       1     |  "18Kb"   |    16384    |    14-bit    |    1-bit   --
   -----------------------------------------------------------------------


   BRAM_SDP_MACRO_inst : BRAM_SDP_MACRO
   generic map (
      BRAM_SIZE => "18Kb", -- Target BRAM, "18Kb" or "36Kb" 
      DEVICE => "7SERIES", -- Target device: "VIRTEX5", "VIRTEX6", "7SERIES", "SPARTAN6" 
      WRITE_WIDTH => 23,    -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
      READ_WIDTH => 23,     -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
      DO_REG => 1, -- Optional output register (0 or 1)
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY", 
                                    -- "GENERATE_X_ONLY" or "NONE"       
      SRVAL => X"101010101010101010", --  Set/Reset value for port output
      WRITE_MODE => "READ_FIRST", -- Specify "READ_FIRST" for same clock or synchronous clocks
                                   --  Specify "WRITE_FIRST for asynchrononous clocks on ports
      INIT => X"000000000000000000", --  Initial values on output port
      -- The following INIT_xx declarations specify the initial contents of the RAM
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      
      -- The next set of INIT_xx are valid when configured as 36Kb
      INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
      
      -- The next set of INITP_xx are for the parity bits
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      
      -- The next set of INIT_xx are valid when configured as 36Kb
      INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO => q,         -- Output read data port, width defined by READ_WIDTH parameter
      DI => d.data,         -- Input write data port, width defined by WRITE_WIDTH parameter
      RDADDR => d.raddr, -- Input read address, width defined by read port depth
      RDCLK => clk,   -- 1-bit input read clock
      RDEN => d.ren,     -- 1-bit input read port enable
      REGCE => '1',   -- 1-bit input read output register enable
      RST => '0',       -- 1-bit input reset 
      WE => d.wen & d.wen & d.wen & d.wen,         -- Input write enable, width defined by write port depth
      WRADDR => d.waddr, -- Input write address, width defined by write port depth
      WRCLK => clk,   -- 1-bit input write clock
      WREN => d.wen      -- 1-bit input write port enable
   );
   -- End of BRAM_SDP_MACRO_inst instantiation
--read: process(clk)
--begin
--    if rising_edge(clk)
--    then
--        if d.ren = '1'
--        then
--            q <= storage(to_integer(unsigned(d.raddr)));
--        else
--            q <= (others => '0');
--        end if;
--    end if;
--end process;

--write: process(clk)
--begin
--    if rising_edge(clk)
--    then
--        if d.wen = '1'
--        then
--            storage(to_integer(unsigned(d.waddr))) <= d.data;
--        end if;
--    end if;
--end process;

--   raddr(13 downto 5) <= d.raddr;
--   raddr(4 downto 0) <= "00000";
--   waddr(13 downto 5) <= d.waddr;
--   waddr(4 downto 0) <= "00000";
--   din(31 downto 23) <= "000000000";
--   din(22 downto 0) <= d.data;
--   q <= dout(22 downto 0);

--   RAMB18E1_inst : RAMB18E1
--   generic map (
--      -- Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
--      RDADDR_COLLISION_HWCONFIG => "PERFORMANCE",
--      -- Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
--      SIM_COLLISION_CHECK => "ALL",
--      -- DOA_REG, DOB_REG: Optional output register (0 or 1)
--      DOA_REG => 1,
--      DOB_REG => 1,
--      -- INITP_00 to INITP_07: Initial contents of parity memory array
--      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      -- INIT_00 to INIT_3F: Initial contents of data memory array
--      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      -- INIT_A, INIT_B: Initial values on output ports
--      INIT_A => X"00000",
--      INIT_B => X"00000",
--      -- Initialization File: RAM initialization file
--      INIT_FILE => "NONE",
--      -- RAM Mode: "SDP" or "TDP" 
--      RAM_MODE => "SDP",
--      -- READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
--      READ_WIDTH_A => 32,                                                              -- 0-72
--      READ_WIDTH_B => 0,                                                               -- 0-18
--      WRITE_WIDTH_A => 0,                                                              -- 0-18
--      WRITE_WIDTH_B => 32,                                                             -- 0-72
--      -- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
--      RSTREG_PRIORITY_A => "REGCE",
--      RSTREG_PRIORITY_B => "REGCE",
--      -- SRVAL_A, SRVAL_B: Set/reset value for output
--      SRVAL_A => X"00000",
--      SRVAL_B => X"00000",
--      -- Simulation Device: Must be set to "7SERIES" for simulation behavior
--      SIM_DEVICE => "7SERIES",
--      -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
--      WRITE_MODE_A => "READ_FIRST",
--      WRITE_MODE_B => "READ_FIRST" 
--   )
--   port map (
--      -- Port A Data: 16-bit (each) output: Port A data
--      DOADO => dout(15 downto 0),     -- 16-bit output: A port data/LSB data
--      DOPADOP => open,                -- 2-bit output: A port parity/LSB parity
--      -- Port B Data: 16-bit (each) output: Port B data
--      DOBDO => dout(31 downto 16),    -- 16-bit output: B port data/MSB data
--      DOPBDOP => open,                -- 2-bit output: B port parity/MSB parity
--      -- Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals (read port
--      -- when RAM_MODE="SDP")
--      ADDRARDADDR => raddr,           -- 14-bit input: A port address/Read address
--      CLKARDCLK => clk,               -- 1-bit input: A port clock/Read clock
--      ENARDEN => d.ren,               -- 1-bit input: A port enable/Read enable
--      REGCEAREGCE => '1',             -- 1-bit input: A port register enable/Register enable
--      RSTRAMARSTRAM => '0',           -- 1-bit input: A port set/reset
--      RSTREGARSTREG => '0',           -- 1-bit input: A port register set/reset
--      WEA => "00",                    -- 2-bit input: A port write enable
--      -- Port A Data: 16-bit (each) input: Port A data
--      DIADI => din(15 downto 0),      -- 16-bit input: A port data/LSB data
--      DIPADIP => "00",                -- 2-bit input: A port parity/LSB parity
--      -- Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals (write port
--      -- when RAM_MODE="SDP")
--      ADDRBWRADDR => waddr,           -- 14-bit input: B port address/Write address
--      CLKBWRCLK => clk,               -- 1-bit input: B port clock/Write clock
--      ENBWREN => d.wen,               -- 1-bit input: B port enable/Write enable
--      REGCEB => '1',                  -- 1-bit input: B port register enable
--      RSTRAMB => '0',                 -- 1-bit input: B port set/reset
--      RSTREGB => '0',                 -- 1-bit input: B port register set/reset
--      WEBWE => (others => d.wen),     -- 4-bit input: B port write enable/Write enable
--      -- Port B Data: 16-bit (each) input: Port B data
--      DIBDI => din(31 downto 16),     -- 16-bit input: B port data/MSB data
--      DIPBDIP => "00"                 -- 2-bit input: B port parity/MSB parity
--   );

end Behavioral;
